// C5G_QSYS.v

// Generated using ACDS version 13.1 162 at 2017.01.01.19:25:14

`timescale 1 ps / 1 ps
module C5G_QSYS (
		input  wire        clk_clk,                                                      //                              clk.clk
		input  wire        reset_reset_n,                                                //                            reset.reset_n
		output wire [9:0]  memory_mem_ca,                                                //                           memory.mem_ca
		output wire [0:0]  memory_mem_ck,                                                //                                 .mem_ck
		output wire [0:0]  memory_mem_ck_n,                                              //                                 .mem_ck_n
		output wire [0:0]  memory_mem_cke,                                               //                                 .mem_cke
		output wire [0:0]  memory_mem_cs_n,                                              //                                 .mem_cs_n
		output wire [3:0]  memory_mem_dm,                                                //                                 .mem_dm
		inout  wire [31:0] memory_mem_dq,                                                //                                 .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                               //                                 .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                             //                                 .mem_dqs_n
		input  wire        oct_rzqin,                                                    //                              oct.rzqin
		output wire        mem_if_lpddr2_emif_status_local_init_done,                    //        mem_if_lpddr2_emif_status.local_init_done
		output wire        mem_if_lpddr2_emif_status_local_cal_success,                  //                                 .local_cal_success
		output wire        mem_if_lpddr2_emif_status_local_cal_fail,                     //                                 .local_cal_fail
		input  wire [3:0]  key_external_connection_export,                               //          key_external_connection.export
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_mem_clk,                   //   mem_if_lpddr2_emif_pll_sharing.pll_mem_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_write_clk,                 //                                 .pll_write_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_locked,                    //                                 .pll_locked
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_write_clk_pre_phy_clk,     //                                 .pll_write_clk_pre_phy_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_addr_cmd_clk,              //                                 .pll_addr_cmd_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_avl_clk,                   //                                 .pll_avl_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_config_clk,                //                                 .pll_config_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_mem_phy_clk,               //                                 .pll_mem_phy_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_afi_phy_clk,                   //                                 .afi_phy_clk
		output wire        mem_if_lpddr2_emif_pll_sharing_pll_avl_phy_clk,               //                                 .pll_avl_phy_clk
		output wire        mem_if_lpddr2_emif_avl_0_waitrequest_n,                       //         mem_if_lpddr2_emif_avl_0.waitrequest_n
		input  wire        mem_if_lpddr2_emif_avl_0_beginbursttransfer,                  //                                 .beginbursttransfer
		input  wire [26:0] mem_if_lpddr2_emif_avl_0_address,                             //                                 .address
		output wire        mem_if_lpddr2_emif_avl_0_readdatavalid,                       //                                 .readdatavalid
		output wire [31:0] mem_if_lpddr2_emif_avl_0_readdata,                            //                                 .readdata
		input  wire [31:0] mem_if_lpddr2_emif_avl_0_writedata,                           //                                 .writedata
		input  wire [3:0]  mem_if_lpddr2_emif_avl_0_byteenable,                          //                                 .byteenable
		input  wire        mem_if_lpddr2_emif_avl_0_read,                                //                                 .read
		input  wire        mem_if_lpddr2_emif_avl_0_write,                               //                                 .write
		input  wire [2:0]  mem_if_lpddr2_emif_avl_0_burstcount,                          //                                 .burstcount
		input  wire        mm_clock_crossing_bridge_0_m0_waitrequest,                    //    mm_clock_crossing_bridge_0_m0.waitrequest
		input  wire [31:0] mm_clock_crossing_bridge_0_m0_readdata,                       //                                 .readdata
		input  wire        mm_clock_crossing_bridge_0_m0_readdatavalid,                  //                                 .readdatavalid
		output wire [3:0]  mm_clock_crossing_bridge_0_m0_burstcount,                     //                                 .burstcount
		output wire [31:0] mm_clock_crossing_bridge_0_m0_writedata,                      //                                 .writedata
		output wire [28:0] mm_clock_crossing_bridge_0_m0_address,                        //                                 .address
		output wire        mm_clock_crossing_bridge_0_m0_write,                          //                                 .write
		output wire        mm_clock_crossing_bridge_0_m0_read,                           //                                 .read
		output wire [3:0]  mm_clock_crossing_bridge_0_m0_byteenable,                     //                                 .byteenable
		output wire        mm_clock_crossing_bridge_0_m0_debugaccess,                    //                                 .debugaccess
		input  wire        uart_usb_rxd,                                                 //                         uart_usb.rxd
		output wire        uart_usb_txd,                                                 //                                 .txd
		output wire [7:0]  led_green_export,                                             //                        led_green.export
		output wire [9:0]  led_red_export,                                               //                          led_red.export
		output wire        sd_card_cs,                                                   //                          sd_card.cs
		output wire        sd_card_sclk,                                                 //                                 .sclk
		output wire        sd_card_mosi,                                                 //                                 .mosi
		input  wire        sd_card_miso,                                                 //                                 .miso
		input  wire        sd_card_cd,                                                   //                                 .cd
		input  wire        sd_card_wp,                                                   //                                 .wp
		inout  wire [15:0] tristate_conduit_bridge_sram_out_sram_tcm_data_out,           // tristate_conduit_bridge_sram_out.sram_tcm_data_out
		output wire [18:0] tristate_conduit_bridge_sram_out_sram_tcm_address_out,        //                                 .sram_tcm_address_out
		output wire [0:0]  tristate_conduit_bridge_sram_out_sram_tcm_outputenable_n_out, //                                 .sram_tcm_outputenable_n_out
		output wire [0:0]  tristate_conduit_bridge_sram_out_sram_tcm_chipselect_n_out,   //                                 .sram_tcm_chipselect_n_out
		output wire [1:0]  tristate_conduit_bridge_sram_out_sram_tcm_byteenable_n_out,   //                                 .sram_tcm_byteenable_n_out
		output wire [0:0]  tristate_conduit_bridge_sram_out_sram_tcm_write_n_out,        //                                 .sram_tcm_write_n_out
		input  wire [9:0]  switches_export                                               //                         switches.export
	);

	wire         mem_if_lpddr2_emif_afi_half_clk_clk;                               // mem_if_lpddr2_emif:afi_half_clk -> [mem_if_lpddr2_emif:mp_cmd_clk_0_clk, mem_if_lpddr2_emif:mp_rfifo_clk_0_clk, mem_if_lpddr2_emif:mp_wfifo_clk_0_clk, mm_clock_crossing_bridge_0:m0_clk, rst_controller_002:clk]
	wire         mem_if_lpddr2_emif_afi_reset_reset;                                // mem_if_lpddr2_emif:afi_reset_n -> [mem_if_lpddr2_emif:mp_cmd_reset_n_0_reset_n, mem_if_lpddr2_emif:mp_rfifo_reset_n_0_reset_n, mem_if_lpddr2_emif:mp_wfifo_reset_n_0_reset_n, rst_controller_002:reset_in0]
	wire         sram_tcm_chipselect_n_out;                                         // sram:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_0:tcs0_chipselect_n_out
	wire         sram_tcm_grant;                                                    // tristate_conduit_pin_sharer_0:tcs0_grant -> sram:tcm_grant
	wire         sram_tcm_data_outen;                                               // sram:tcm_data_outen -> tristate_conduit_pin_sharer_0:tcs0_data_outen
	wire         sram_tcm_outputenable_n_out;                                       // sram:tcm_outputenable_n_out -> tristate_conduit_pin_sharer_0:tcs0_outputenable_n_out
	wire         sram_tcm_request;                                                  // sram:tcm_request -> tristate_conduit_pin_sharer_0:tcs0_request
	wire  [15:0] sram_tcm_data_out;                                                 // sram:tcm_data_out -> tristate_conduit_pin_sharer_0:tcs0_data_out
	wire         sram_tcm_write_n_out;                                              // sram:tcm_write_n_out -> tristate_conduit_pin_sharer_0:tcs0_write_n_out
	wire  [18:0] sram_tcm_address_out;                                              // sram:tcm_address_out -> tristate_conduit_pin_sharer_0:tcs0_address_out
	wire  [15:0] sram_tcm_data_in;                                                  // tristate_conduit_pin_sharer_0:tcs0_data_in -> sram:tcm_data_in
	wire   [1:0] sram_tcm_byteenable_n_out;                                         // sram:tcm_byteenable_n_out -> tristate_conduit_pin_sharer_0:tcs0_byteenable_n_out
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_write_n_out_out;        // tristate_conduit_pin_sharer_0:sram_tcm_write_n_out -> tristate_conduit_bridge_0:tcs_sram_tcm_write_n_out
	wire  [18:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_address_out_out;        // tristate_conduit_pin_sharer_0:sram_tcm_address_out -> tristate_conduit_bridge_0:tcs_sram_tcm_address_out
	wire         tristate_conduit_pin_sharer_0_tcm_grant;                           // tristate_conduit_bridge_0:grant -> tristate_conduit_pin_sharer_0:grant
	wire         tristate_conduit_pin_sharer_0_tcm_request;                         // tristate_conduit_pin_sharer_0:request -> tristate_conduit_bridge_0:request
	wire   [1:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_byteenable_n_out_out;   // tristate_conduit_pin_sharer_0:sram_tcm_byteenable_n_out -> tristate_conduit_bridge_0:tcs_sram_tcm_byteenable_n_out
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_outputenable_n_out_out; // tristate_conduit_pin_sharer_0:sram_tcm_outputenable_n_out -> tristate_conduit_bridge_0:tcs_sram_tcm_outputenable_n_out
	wire         tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_outen;         // tristate_conduit_pin_sharer_0:sram_tcm_data_outen -> tristate_conduit_bridge_0:tcs_sram_tcm_data_outen
	wire  [15:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_in;            // tristate_conduit_bridge_0:tcs_sram_tcm_data_in -> tristate_conduit_pin_sharer_0:sram_tcm_data_in
	wire  [15:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_out;           // tristate_conduit_pin_sharer_0:sram_tcm_data_out -> tristate_conduit_bridge_0:tcs_sram_tcm_data_out
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_sram_tcm_chipselect_n_out_out;   // tristate_conduit_pin_sharer_0:sram_tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_sram_tcm_chipselect_n_out
	wire  [15:0] mm_interconnect_0_uart_usb_s1_writedata;                           // mm_interconnect_0:uart_usb_s1_writedata -> uart_usb:writedata
	wire   [2:0] mm_interconnect_0_uart_usb_s1_address;                             // mm_interconnect_0:uart_usb_s1_address -> uart_usb:address
	wire         mm_interconnect_0_uart_usb_s1_chipselect;                          // mm_interconnect_0:uart_usb_s1_chipselect -> uart_usb:chipselect
	wire         mm_interconnect_0_uart_usb_s1_write;                               // mm_interconnect_0:uart_usb_s1_write -> uart_usb:write_n
	wire         mm_interconnect_0_uart_usb_s1_read;                                // mm_interconnect_0:uart_usb_s1_read -> uart_usb:read_n
	wire  [15:0] mm_interconnect_0_uart_usb_s1_readdata;                            // uart_usb:readdata -> mm_interconnect_0:uart_usb_s1_readdata
	wire         mm_interconnect_0_uart_usb_s1_begintransfer;                       // mm_interconnect_0:uart_usb_s1_begintransfer -> uart_usb:begintransfer
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                     // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                       // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                         // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_onchip_memory2_s1_write;                         // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                      // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         nios2_qsys_data_master_waitrequest;                                // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                                  // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [30:0] nios2_qsys_data_master_address;                                    // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire         nios2_qsys_data_master_write;                                      // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire         nios2_qsys_data_master_read;                                       // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire  [31:0] nios2_qsys_data_master_readdata;                                   // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                                // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                              // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                                 // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;                // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;                  // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;               // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire         mm_interconnect_0_epcs_epcs_control_port_write;                    // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire         mm_interconnect_0_epcs_epcs_control_port_read;                     // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;                 // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;               // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire  [31:0] mm_interconnect_0_led_green_s1_writedata;                          // mm_interconnect_0:led_green_s1_writedata -> led_green:writedata
	wire   [1:0] mm_interconnect_0_led_green_s1_address;                            // mm_interconnect_0:led_green_s1_address -> led_green:address
	wire         mm_interconnect_0_led_green_s1_chipselect;                         // mm_interconnect_0:led_green_s1_chipselect -> led_green:chipselect
	wire         mm_interconnect_0_led_green_s1_write;                              // mm_interconnect_0:led_green_s1_write -> led_green:write_n
	wire  [31:0] mm_interconnect_0_led_green_s1_readdata;                           // led_green:readdata -> mm_interconnect_0:led_green_s1_readdata
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                                // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                  // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_key_s1_chipselect;                               // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire         mm_interconnect_0_key_s1_write;                                    // mm_interconnect_0:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                 // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest;        // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;          // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;            // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_write;              // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_read;               // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;           // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess;        // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;         // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire   [1:0] mm_interconnect_0_switches_s1_address;                             // mm_interconnect_0:switches_s1_address -> switches:address
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                            // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_spi_master_0_s1_writedata;                       // mm_interconnect_0:spi_master_0_s1_writedata -> spi_master_0:writedata
	wire   [2:0] mm_interconnect_0_spi_master_0_s1_address;                         // mm_interconnect_0:spi_master_0_s1_address -> spi_master_0:address
	wire         mm_interconnect_0_spi_master_0_s1_chipselect;                      // mm_interconnect_0:spi_master_0_s1_chipselect -> spi_master_0:chipselect
	wire         mm_interconnect_0_spi_master_0_s1_write;                           // mm_interconnect_0:spi_master_0_s1_write -> spi_master_0:write
	wire         mm_interconnect_0_spi_master_0_s1_read;                            // mm_interconnect_0:spi_master_0_s1_read -> spi_master_0:read
	wire  [31:0] mm_interconnect_0_spi_master_0_s1_readdata;                        // spi_master_0:readdata -> mm_interconnect_0:spi_master_0_s1_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [30:0] nios2_qsys_instruction_master_address;                             // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                                // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                            // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire  [31:0] mm_interconnect_0_led_red_s1_writedata;                            // mm_interconnect_0:led_red_s1_writedata -> led_red:writedata
	wire   [1:0] mm_interconnect_0_led_red_s1_address;                              // mm_interconnect_0:led_red_s1_address -> led_red:address
	wire         mm_interconnect_0_led_red_s1_chipselect;                           // mm_interconnect_0:led_red_s1_chipselect -> led_red:chipselect
	wire         mm_interconnect_0_led_red_s1_write;                                // mm_interconnect_0:led_red_s1_write -> led_red:write_n
	wire  [31:0] mm_interconnect_0_led_red_s1_readdata;                             // led_red:readdata -> mm_interconnect_0:led_red_s1_readdata
	wire         mm_interconnect_0_sram_uas_waitrequest;                            // sram:uas_waitrequest -> mm_interconnect_0:sram_uas_waitrequest
	wire   [1:0] mm_interconnect_0_sram_uas_burstcount;                             // mm_interconnect_0:sram_uas_burstcount -> sram:uas_burstcount
	wire  [15:0] mm_interconnect_0_sram_uas_writedata;                              // mm_interconnect_0:sram_uas_writedata -> sram:uas_writedata
	wire  [18:0] mm_interconnect_0_sram_uas_address;                                // mm_interconnect_0:sram_uas_address -> sram:uas_address
	wire         mm_interconnect_0_sram_uas_lock;                                   // mm_interconnect_0:sram_uas_lock -> sram:uas_lock
	wire         mm_interconnect_0_sram_uas_write;                                  // mm_interconnect_0:sram_uas_write -> sram:uas_write
	wire         mm_interconnect_0_sram_uas_read;                                   // mm_interconnect_0:sram_uas_read -> sram:uas_read
	wire  [15:0] mm_interconnect_0_sram_uas_readdata;                               // sram:uas_readdata -> mm_interconnect_0:sram_uas_readdata
	wire         mm_interconnect_0_sram_uas_debugaccess;                            // mm_interconnect_0:sram_uas_debugaccess -> sram:uas_debugaccess
	wire         mm_interconnect_0_sram_uas_readdatavalid;                          // sram:uas_readdatavalid -> mm_interconnect_0:sram_uas_readdatavalid
	wire   [1:0] mm_interconnect_0_sram_uas_byteenable;                             // mm_interconnect_0:sram_uas_byteenable -> sram:uas_byteenable
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                              // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                             // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                                  // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                               // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest;       // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount;        // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata;         // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire  [28:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address;           // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write;             // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read;              // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata;          // mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess;       // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid;     // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable;        // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire         irq_mapper_receiver0_irq;                                          // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                          // key:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                          // uart_usb:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                          // epcs:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                              // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [nios2_qsys:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_jtag_debug_module_reset_reset;                          // nios2_qsys:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [epcs:reset_n, jtag_uart:rst_n, key:reset_n, led_green:reset_n, led_red:reset_n, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:onchip_memory2_reset1_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator_001:in_reset, spi_master_0:reset, sram:reset_reset, switches:reset_n, sysid_qsys:reset_n, timer:reset_n, tristate_conduit_bridge_0:reset, tristate_conduit_pin_sharer_0:reset_reset, uart_usb:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                            // rst_controller_001:reset_req -> [epcs:reset_req, onchip_memory2:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> mm_clock_crossing_bridge_0:m0_reset

	C5G_QSYS_nios2_qsys nios2_qsys (
		.clk                                   (clk_clk),                                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	C5G_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	C5G_QSYS_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	C5G_QSYS_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	C5G_QSYS_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	C5G_QSYS_mem_if_lpddr2_emif mem_if_lpddr2_emif (
		.pll_ref_clk                (clk_clk),                                                  //        pll_ref_clk.clk
		.global_reset_n             (reset_reset_n),                                            //       global_reset.reset_n
		.soft_reset_n               (reset_reset_n),                                            //         soft_reset.reset_n
		.afi_clk                    (),                                                         //            afi_clk.clk
		.afi_half_clk               (mem_if_lpddr2_emif_afi_half_clk_clk),                      //       afi_half_clk.clk
		.afi_reset_n                (mem_if_lpddr2_emif_afi_reset_reset),                       //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                         //   afi_reset_export.reset_n
		.mem_ca                     (memory_mem_ca),                                            //             memory.mem_ca
		.mem_ck                     (memory_mem_ck),                                            //                   .mem_ck
		.mem_ck_n                   (memory_mem_ck_n),                                          //                   .mem_ck_n
		.mem_cke                    (memory_mem_cke),                                           //                   .mem_cke
		.mem_cs_n                   (memory_mem_cs_n),                                          //                   .mem_cs_n
		.mem_dm                     (memory_mem_dm),                                            //                   .mem_dm
		.mem_dq                     (memory_mem_dq),                                            //                   .mem_dq
		.mem_dqs                    (memory_mem_dqs),                                           //                   .mem_dqs
		.mem_dqs_n                  (memory_mem_dqs_n),                                         //                   .mem_dqs_n
		.avl_ready_0                (mem_if_lpddr2_emif_avl_0_waitrequest_n),                   //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mem_if_lpddr2_emif_avl_0_beginbursttransfer),              //                   .beginbursttransfer
		.avl_addr_0                 (mem_if_lpddr2_emif_avl_0_address),                         //                   .address
		.avl_rdata_valid_0          (mem_if_lpddr2_emif_avl_0_readdatavalid),                   //                   .readdatavalid
		.avl_rdata_0                (mem_if_lpddr2_emif_avl_0_readdata),                        //                   .readdata
		.avl_wdata_0                (mem_if_lpddr2_emif_avl_0_writedata),                       //                   .writedata
		.avl_be_0                   (mem_if_lpddr2_emif_avl_0_byteenable),                      //                   .byteenable
		.avl_read_req_0             (mem_if_lpddr2_emif_avl_0_read),                            //                   .read
		.avl_write_req_0            (mem_if_lpddr2_emif_avl_0_write),                           //                   .write
		.avl_size_0                 (mem_if_lpddr2_emif_avl_0_burstcount),                      //                   .burstcount
		.mp_cmd_clk_0_clk           (mem_if_lpddr2_emif_afi_half_clk_clk),                      //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (mem_if_lpddr2_emif_afi_reset_reset),                       //   mp_cmd_reset_n_0.reset_n
		.mp_rfifo_clk_0_clk         (mem_if_lpddr2_emif_afi_half_clk_clk),                      //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (mem_if_lpddr2_emif_afi_reset_reset),                       // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (mem_if_lpddr2_emif_afi_half_clk_clk),                      //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (mem_if_lpddr2_emif_afi_reset_reset),                       // mp_wfifo_reset_n_0.reset_n
		.local_init_done            (mem_if_lpddr2_emif_status_local_init_done),                //             status.local_init_done
		.local_cal_success          (mem_if_lpddr2_emif_status_local_cal_success),              //                   .local_cal_success
		.local_cal_fail             (mem_if_lpddr2_emif_status_local_cal_fail),                 //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                                //                oct.rzqin
		.pll_mem_clk                (mem_if_lpddr2_emif_pll_sharing_pll_mem_clk),               //        pll_sharing.pll_mem_clk
		.pll_write_clk              (mem_if_lpddr2_emif_pll_sharing_pll_write_clk),             //                   .pll_write_clk
		.pll_locked                 (mem_if_lpddr2_emif_pll_sharing_pll_locked),                //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (mem_if_lpddr2_emif_pll_sharing_pll_write_clk_pre_phy_clk), //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (mem_if_lpddr2_emif_pll_sharing_pll_addr_cmd_clk),          //                   .pll_addr_cmd_clk
		.pll_avl_clk                (mem_if_lpddr2_emif_pll_sharing_pll_avl_clk),               //                   .pll_avl_clk
		.pll_config_clk             (mem_if_lpddr2_emif_pll_sharing_pll_config_clk),            //                   .pll_config_clk
		.pll_mem_phy_clk            (mem_if_lpddr2_emif_pll_sharing_pll_mem_phy_clk),           //                   .pll_mem_phy_clk
		.afi_phy_clk                (mem_if_lpddr2_emif_pll_sharing_afi_phy_clk),               //                   .afi_phy_clk
		.pll_avl_phy_clk            (mem_if_lpddr2_emif_pll_sharing_pll_avl_phy_clk)            //                   .pll_avl_phy_clk
	);

	C5G_QSYS_key key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (29),
		.BURSTCOUNT_WIDTH    (4),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (mem_if_lpddr2_emif_afi_half_clk_clk),                           //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (clk_clk),                                                       //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	C5G_QSYS_uart_usb uart_usb (
		.clk           (clk_clk),                                     //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_usb_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_usb_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_usb_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_usb_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_usb_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_usb_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_usb_s1_readdata),      //                    .readdata
		.dataavailable (),                                            //                    .dataavailable
		.readyfordata  (),                                            //                    .readyfordata
		.rxd           (uart_usb_rxd),                                // external_connection.export
		.txd           (uart_usb_txd),                                //                    .export
		.irq           (irq_mapper_receiver3_irq)                     //                 irq.irq
	);

	C5G_QSYS_led_green led_green (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_green_s1_readdata),   //                    .readdata
		.out_port   (led_green_export)                           // external_connection.export
	);

	C5G_QSYS_led_red led_red (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_red_s1_readdata),   //                    .readdata
		.out_port   (led_red_export)                           // external_connection.export
	);

	spi_master_if spi_master_0 (
		.reset      (rst_controller_001_reset_out_reset),           //    reset.reset
		.clk        (clk_clk),                                      //      clk.clk
		.chipselect (mm_interconnect_0_spi_master_0_s1_chipselect), //       s1.chipselect
		.address    (mm_interconnect_0_spi_master_0_s1_address),    //         .address
		.write      (mm_interconnect_0_spi_master_0_s1_write),      //         .write
		.writedata  (mm_interconnect_0_spi_master_0_s1_writedata),  //         .writedata
		.read       (mm_interconnect_0_spi_master_0_s1_read),       //         .read
		.readdata   (mm_interconnect_0_spi_master_0_s1_readdata),   //         .readdata
		.cs         (sd_card_cs),                                   // external.export
		.sclk       (sd_card_sclk),                                 //         .export
		.mosi       (sd_card_mosi),                                 //         .export
		.miso       (sd_card_miso),                                 //         .export
		.cd         (sd_card_cd),                                   //         .export
		.wp         (sd_card_wp)                                    //         .export
	);

	C5G_QSYS_sram #(
		.TCM_ADDRESS_W                  (19),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (10),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (10),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram (
		.clk_clk                (clk_clk),                                  //   clk.clk
		.reset_reset            (rst_controller_001_reset_out_reset),       // reset.reset
		.uas_address            (mm_interconnect_0_sram_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_0_sram_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_0_sram_uas_read),          //      .read
		.uas_write              (mm_interconnect_0_sram_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_0_sram_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_0_sram_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_0_sram_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_0_sram_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_0_sram_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_0_sram_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_0_sram_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (sram_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (sram_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (sram_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request            (sram_tcm_request),                         //      .request
		.tcm_grant              (sram_tcm_grant),                           //      .grant
		.tcm_address_out        (sram_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out   (sram_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out           (sram_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (sram_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (sram_tcm_data_in)                          //      .data_in
	);

	C5G_QSYS_tristate_conduit_pin_sharer_0 tristate_conduit_pin_sharer_0 (
		.clk_clk                     (clk_clk),                                                           //   clk.clk
		.reset_reset                 (rst_controller_001_reset_out_reset),                                // reset.reset
		.request                     (tristate_conduit_pin_sharer_0_tcm_request),                         //   tcm.request
		.grant                       (tristate_conduit_pin_sharer_0_tcm_grant),                           //      .grant
		.sram_tcm_address_out        (tristate_conduit_pin_sharer_0_tcm_sram_tcm_address_out_out),        //      .sram_tcm_address_out_out
		.sram_tcm_outputenable_n_out (tristate_conduit_pin_sharer_0_tcm_sram_tcm_outputenable_n_out_out), //      .sram_tcm_outputenable_n_out_out
		.sram_tcm_byteenable_n_out   (tristate_conduit_pin_sharer_0_tcm_sram_tcm_byteenable_n_out_out),   //      .sram_tcm_byteenable_n_out_out
		.sram_tcm_write_n_out        (tristate_conduit_pin_sharer_0_tcm_sram_tcm_write_n_out_out),        //      .sram_tcm_write_n_out_out
		.sram_tcm_data_out           (tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_out),           //      .sram_tcm_data_out_out
		.sram_tcm_data_in            (tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_in),            //      .sram_tcm_data_out_in
		.sram_tcm_data_outen         (tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_outen),         //      .sram_tcm_data_out_outen
		.sram_tcm_chipselect_n_out   (tristate_conduit_pin_sharer_0_tcm_sram_tcm_chipselect_n_out_out),   //      .sram_tcm_chipselect_n_out_out
		.tcs0_request                (sram_tcm_request),                                                  //  tcs0.request
		.tcs0_grant                  (sram_tcm_grant),                                                    //      .grant
		.tcs0_address_out            (sram_tcm_address_out),                                              //      .address_out
		.tcs0_outputenable_n_out     (sram_tcm_outputenable_n_out),                                       //      .outputenable_n_out
		.tcs0_byteenable_n_out       (sram_tcm_byteenable_n_out),                                         //      .byteenable_n_out
		.tcs0_write_n_out            (sram_tcm_write_n_out),                                              //      .write_n_out
		.tcs0_data_out               (sram_tcm_data_out),                                                 //      .data_out
		.tcs0_data_in                (sram_tcm_data_in),                                                  //      .data_in
		.tcs0_data_outen             (sram_tcm_data_outen),                                               //      .data_outen
		.tcs0_chipselect_n_out       (sram_tcm_chipselect_n_out)                                          //      .chipselect_n_out
	);

	C5G_QSYS_tristate_conduit_bridge_0 tristate_conduit_bridge_0 (
		.clk                             (clk_clk),                                                           //   clk.clk
		.reset                           (rst_controller_001_reset_out_reset),                                // reset.reset
		.request                         (tristate_conduit_pin_sharer_0_tcm_request),                         //   tcs.request
		.grant                           (tristate_conduit_pin_sharer_0_tcm_grant),                           //      .grant
		.tcs_sram_tcm_data_out           (tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_out),           //      .sram_tcm_data_out_out
		.tcs_sram_tcm_data_outen         (tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_outen),         //      .sram_tcm_data_out_outen
		.tcs_sram_tcm_data_in            (tristate_conduit_pin_sharer_0_tcm_sram_tcm_data_out_in),            //      .sram_tcm_data_out_in
		.tcs_sram_tcm_address_out        (tristate_conduit_pin_sharer_0_tcm_sram_tcm_address_out_out),        //      .sram_tcm_address_out_out
		.tcs_sram_tcm_outputenable_n_out (tristate_conduit_pin_sharer_0_tcm_sram_tcm_outputenable_n_out_out), //      .sram_tcm_outputenable_n_out_out
		.tcs_sram_tcm_chipselect_n_out   (tristate_conduit_pin_sharer_0_tcm_sram_tcm_chipselect_n_out_out),   //      .sram_tcm_chipselect_n_out_out
		.tcs_sram_tcm_byteenable_n_out   (tristate_conduit_pin_sharer_0_tcm_sram_tcm_byteenable_n_out_out),   //      .sram_tcm_byteenable_n_out_out
		.tcs_sram_tcm_write_n_out        (tristate_conduit_pin_sharer_0_tcm_sram_tcm_write_n_out_out),        //      .sram_tcm_write_n_out_out
		.sram_tcm_data_out               (tristate_conduit_bridge_sram_out_sram_tcm_data_out),                //   out.sram_tcm_data_out
		.sram_tcm_address_out            (tristate_conduit_bridge_sram_out_sram_tcm_address_out),             //      .sram_tcm_address_out
		.sram_tcm_outputenable_n_out     (tristate_conduit_bridge_sram_out_sram_tcm_outputenable_n_out),      //      .sram_tcm_outputenable_n_out
		.sram_tcm_chipselect_n_out       (tristate_conduit_bridge_sram_out_sram_tcm_chipselect_n_out),        //      .sram_tcm_chipselect_n_out
		.sram_tcm_byteenable_n_out       (tristate_conduit_bridge_sram_out_sram_tcm_byteenable_n_out),        //      .sram_tcm_byteenable_n_out
		.sram_tcm_write_n_out            (tristate_conduit_bridge_sram_out_sram_tcm_write_n_out)              //      .sram_tcm_write_n_out
	);

	C5G_QSYS_epcs epcs (
		.clk           (clk_clk),                                             //               clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                 //             reset.reset_n
		.reset_req     (rst_controller_001_reset_out_reset_req),              //                  .reset_req
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver4_irq)                             //               irq.irq
	);

	C5G_QSYS_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	C5G_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_125_clk_clk                                   (clk_clk),                                                       //                                 clk_125_clk.clk
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                                //    nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.onchip_memory2_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // onchip_memory2_reset1_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                    (nios2_qsys_data_master_address),                                //                      nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest                (nios2_qsys_data_master_waitrequest),                            //                                            .waitrequest
		.nios2_qsys_data_master_byteenable                 (nios2_qsys_data_master_byteenable),                             //                                            .byteenable
		.nios2_qsys_data_master_read                       (nios2_qsys_data_master_read),                                   //                                            .read
		.nios2_qsys_data_master_readdata                   (nios2_qsys_data_master_readdata),                               //                                            .readdata
		.nios2_qsys_data_master_readdatavalid              (nios2_qsys_data_master_readdatavalid),                          //                                            .readdatavalid
		.nios2_qsys_data_master_write                      (nios2_qsys_data_master_write),                                  //                                            .write
		.nios2_qsys_data_master_writedata                  (nios2_qsys_data_master_writedata),                              //                                            .writedata
		.nios2_qsys_data_master_debugaccess                (nios2_qsys_data_master_debugaccess),                            //                                            .debugaccess
		.nios2_qsys_instruction_master_address             (nios2_qsys_instruction_master_address),                         //               nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest         (nios2_qsys_instruction_master_waitrequest),                     //                                            .waitrequest
		.nios2_qsys_instruction_master_read                (nios2_qsys_instruction_master_read),                            //                                            .read
		.nios2_qsys_instruction_master_readdata            (nios2_qsys_instruction_master_readdata),                        //                                            .readdata
		.nios2_qsys_instruction_master_readdatavalid       (nios2_qsys_instruction_master_readdatavalid),                   //                                            .readdatavalid
		.epcs_epcs_control_port_address                    (mm_interconnect_0_epcs_epcs_control_port_address),              //                      epcs_epcs_control_port.address
		.epcs_epcs_control_port_write                      (mm_interconnect_0_epcs_epcs_control_port_write),                //                                            .write
		.epcs_epcs_control_port_read                       (mm_interconnect_0_epcs_epcs_control_port_read),                 //                                            .read
		.epcs_epcs_control_port_readdata                   (mm_interconnect_0_epcs_epcs_control_port_readdata),             //                                            .readdata
		.epcs_epcs_control_port_writedata                  (mm_interconnect_0_epcs_epcs_control_port_writedata),            //                                            .writedata
		.epcs_epcs_control_port_chipselect                 (mm_interconnect_0_epcs_epcs_control_port_chipselect),           //                                            .chipselect
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                 jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                            .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                            .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                            .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                            .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                            .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                            .chipselect
		.key_s1_address                                    (mm_interconnect_0_key_s1_address),                              //                                      key_s1.address
		.key_s1_write                                      (mm_interconnect_0_key_s1_write),                                //                                            .write
		.key_s1_readdata                                   (mm_interconnect_0_key_s1_readdata),                             //                                            .readdata
		.key_s1_writedata                                  (mm_interconnect_0_key_s1_writedata),                            //                                            .writedata
		.key_s1_chipselect                                 (mm_interconnect_0_key_s1_chipselect),                           //                                            .chipselect
		.led_green_s1_address                              (mm_interconnect_0_led_green_s1_address),                        //                                led_green_s1.address
		.led_green_s1_write                                (mm_interconnect_0_led_green_s1_write),                          //                                            .write
		.led_green_s1_readdata                             (mm_interconnect_0_led_green_s1_readdata),                       //                                            .readdata
		.led_green_s1_writedata                            (mm_interconnect_0_led_green_s1_writedata),                      //                                            .writedata
		.led_green_s1_chipselect                           (mm_interconnect_0_led_green_s1_chipselect),                     //                                            .chipselect
		.led_red_s1_address                                (mm_interconnect_0_led_red_s1_address),                          //                                  led_red_s1.address
		.led_red_s1_write                                  (mm_interconnect_0_led_red_s1_write),                            //                                            .write
		.led_red_s1_readdata                               (mm_interconnect_0_led_red_s1_readdata),                         //                                            .readdata
		.led_red_s1_writedata                              (mm_interconnect_0_led_red_s1_writedata),                        //                                            .writedata
		.led_red_s1_chipselect                             (mm_interconnect_0_led_red_s1_chipselect),                       //                                            .chipselect
		.mm_clock_crossing_bridge_0_s0_address             (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //               mm_clock_crossing_bridge_0_s0.address
		.mm_clock_crossing_bridge_0_s0_write               (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //                                            .write
		.mm_clock_crossing_bridge_0_s0_read                (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //                                            .read
		.mm_clock_crossing_bridge_0_s0_readdata            (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //                                            .readdata
		.mm_clock_crossing_bridge_0_s0_writedata           (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //                                            .writedata
		.mm_clock_crossing_bridge_0_s0_burstcount          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //                                            .burstcount
		.mm_clock_crossing_bridge_0_s0_byteenable          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //                                            .byteenable
		.mm_clock_crossing_bridge_0_s0_readdatavalid       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //                                            .readdatavalid
		.mm_clock_crossing_bridge_0_s0_waitrequest         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //                                            .waitrequest
		.mm_clock_crossing_bridge_0_s0_debugaccess         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //                                            .debugaccess
		.nios2_qsys_jtag_debug_module_address              (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),        //                nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write                (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),          //                                            .write
		.nios2_qsys_jtag_debug_module_read                 (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),           //                                            .read
		.nios2_qsys_jtag_debug_module_readdata             (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),       //                                            .readdata
		.nios2_qsys_jtag_debug_module_writedata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),      //                                            .writedata
		.nios2_qsys_jtag_debug_module_byteenable           (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),     //                                            .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest          (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest),    //                                            .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess          (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess),    //                                            .debugaccess
		.onchip_memory2_s1_address                         (mm_interconnect_0_onchip_memory2_s1_address),                   //                           onchip_memory2_s1.address
		.onchip_memory2_s1_write                           (mm_interconnect_0_onchip_memory2_s1_write),                     //                                            .write
		.onchip_memory2_s1_readdata                        (mm_interconnect_0_onchip_memory2_s1_readdata),                  //                                            .readdata
		.onchip_memory2_s1_writedata                       (mm_interconnect_0_onchip_memory2_s1_writedata),                 //                                            .writedata
		.onchip_memory2_s1_byteenable                      (mm_interconnect_0_onchip_memory2_s1_byteenable),                //                                            .byteenable
		.onchip_memory2_s1_chipselect                      (mm_interconnect_0_onchip_memory2_s1_chipselect),                //                                            .chipselect
		.onchip_memory2_s1_clken                           (mm_interconnect_0_onchip_memory2_s1_clken),                     //                                            .clken
		.spi_master_0_s1_address                           (mm_interconnect_0_spi_master_0_s1_address),                     //                             spi_master_0_s1.address
		.spi_master_0_s1_write                             (mm_interconnect_0_spi_master_0_s1_write),                       //                                            .write
		.spi_master_0_s1_read                              (mm_interconnect_0_spi_master_0_s1_read),                        //                                            .read
		.spi_master_0_s1_readdata                          (mm_interconnect_0_spi_master_0_s1_readdata),                    //                                            .readdata
		.spi_master_0_s1_writedata                         (mm_interconnect_0_spi_master_0_s1_writedata),                   //                                            .writedata
		.spi_master_0_s1_chipselect                        (mm_interconnect_0_spi_master_0_s1_chipselect),                  //                                            .chipselect
		.sram_uas_address                                  (mm_interconnect_0_sram_uas_address),                            //                                    sram_uas.address
		.sram_uas_write                                    (mm_interconnect_0_sram_uas_write),                              //                                            .write
		.sram_uas_read                                     (mm_interconnect_0_sram_uas_read),                               //                                            .read
		.sram_uas_readdata                                 (mm_interconnect_0_sram_uas_readdata),                           //                                            .readdata
		.sram_uas_writedata                                (mm_interconnect_0_sram_uas_writedata),                          //                                            .writedata
		.sram_uas_burstcount                               (mm_interconnect_0_sram_uas_burstcount),                         //                                            .burstcount
		.sram_uas_byteenable                               (mm_interconnect_0_sram_uas_byteenable),                         //                                            .byteenable
		.sram_uas_readdatavalid                            (mm_interconnect_0_sram_uas_readdatavalid),                      //                                            .readdatavalid
		.sram_uas_waitrequest                              (mm_interconnect_0_sram_uas_waitrequest),                        //                                            .waitrequest
		.sram_uas_lock                                     (mm_interconnect_0_sram_uas_lock),                               //                                            .lock
		.sram_uas_debugaccess                              (mm_interconnect_0_sram_uas_debugaccess),                        //                                            .debugaccess
		.switches_s1_address                               (mm_interconnect_0_switches_s1_address),                         //                                 switches_s1.address
		.switches_s1_readdata                              (mm_interconnect_0_switches_s1_readdata),                        //                                            .readdata
		.sysid_qsys_control_slave_address                  (mm_interconnect_0_sysid_qsys_control_slave_address),            //                    sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                 (mm_interconnect_0_sysid_qsys_control_slave_readdata),           //                                            .readdata
		.timer_s1_address                                  (mm_interconnect_0_timer_s1_address),                            //                                    timer_s1.address
		.timer_s1_write                                    (mm_interconnect_0_timer_s1_write),                              //                                            .write
		.timer_s1_readdata                                 (mm_interconnect_0_timer_s1_readdata),                           //                                            .readdata
		.timer_s1_writedata                                (mm_interconnect_0_timer_s1_writedata),                          //                                            .writedata
		.timer_s1_chipselect                               (mm_interconnect_0_timer_s1_chipselect),                         //                                            .chipselect
		.uart_usb_s1_address                               (mm_interconnect_0_uart_usb_s1_address),                         //                                 uart_usb_s1.address
		.uart_usb_s1_write                                 (mm_interconnect_0_uart_usb_s1_write),                           //                                            .write
		.uart_usb_s1_read                                  (mm_interconnect_0_uart_usb_s1_read),                            //                                            .read
		.uart_usb_s1_readdata                              (mm_interconnect_0_uart_usb_s1_readdata),                        //                                            .readdata
		.uart_usb_s1_writedata                             (mm_interconnect_0_uart_usb_s1_writedata),                       //                                            .writedata
		.uart_usb_s1_begintransfer                         (mm_interconnect_0_uart_usb_s1_begintransfer),                   //                                            .begintransfer
		.uart_usb_s1_chipselect                            (mm_interconnect_0_uart_usb_s1_chipselect)                       //                                            .chipselect
	);

	C5G_QSYS_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~mem_if_lpddr2_emif_afi_reset_reset), // reset_in0.reset
		.clk            (mem_if_lpddr2_emif_afi_half_clk_clk), //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
